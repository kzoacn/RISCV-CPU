module station(
		input wire clk,	
		output reg busy,
		output reg[6:0] opcode,
		output reg[2:0] fun3,
		output reg[6:0] fun7,
		output reg[31:0] vj,
		output reg[31:0] vk,
		output reg[4:0] qj,
		output reg[4:0] qk,
		output reg[31:0] A
	);


	
endmodule

