module RSREG
